** Profile: "SCHEMATIC1-test"  [ C:\USERS\M R\DESKTOP\AZ MADAR ELEC\s10\pish6\pish6-SCHEMATIC1-test.sim ] 

** Creating circuit file "pish6-SCHEMATIC1-test.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 100ms 0 100u 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\pish6-SCHEMATIC1.net" 


.END
