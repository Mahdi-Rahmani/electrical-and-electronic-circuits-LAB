** Profile: "SCHEMATIC1-tes2"  [ C:\USERS\M R\DESKTOP\AZ MADAR ELEC\s09\az1\az1-SCHEMATIC1-tes2.sim ] 

** Creating circuit file "az1-SCHEMATIC1-tes2.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\az1-SCHEMATIC1.net" 


.END
