** Profile: "SCHEMATIC1-test1"  [ C:\USERS\M R\DESKTOP\AZ MADAR ELEC\elec project\q2\part2-SCHEMATIC1-test1.sim ] 

** Creating circuit file "part2-SCHEMATIC1-test1.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 10000 1u 100k
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\part2-SCHEMATIC1.net" 


.END
