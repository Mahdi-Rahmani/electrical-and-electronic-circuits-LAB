** Profile: "SCHEMATIC1-q1_pishgozarsh2"  [ C:\Users\M R\Desktop\az madar elec\pishgozaresh\q1\pishgozaresh1-SCHEMATIC1-q1_pishgozarsh2.sim ] 

** Creating circuit file "pishgozaresh1-SCHEMATIC1-q1_pishgozarsh2.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1000ns 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\pishgozaresh1-SCHEMATIC1.net" 


.END
