** Profile: "SCHEMATIC1-sim"  [ C:\USERS\M R\DESKTOP\az madar elec\s07\pishGozaresh2\q2-SCHEMATIC1-sim.sim ] 

** Creating circuit file "q2-SCHEMATIC1-sim.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 1000 0.1 200k
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\q2-SCHEMATIC1.net" 


.END
