** Profile: "SCHEMATIC1-q2-1"  [ C:\Users\M R\Desktop\az madar elec\pishgozaresh\q2_2\q2_pishgozaresh-SCHEMATIC1-q2-1.sim ] 

** Creating circuit file "q2_pishgozaresh-SCHEMATIC1-q2-1.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\q2_pishgozaresh-SCHEMATIC1.net" 


.END
