** Profile: "SCHEMATIC1-test"  [ C:\Users\M R\Desktop\az madar elec\s03\pish gozaresh 3\q6-SCHEMATIC1-test.sim ] 

** Creating circuit file "q6-SCHEMATIC1-test.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN PARAM a 1 1k 5 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\q6-SCHEMATIC1.net" 


.END
