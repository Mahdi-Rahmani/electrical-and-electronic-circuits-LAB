** Profile: "SCHEMATIC1-test"  [ C:\USERS\M R\DESKTOP\AZ MADAR ELEC\ELEC PROJECT\q6\IN\part6_2-SCHEMATIC1-test.sim ] 

** Creating circuit file "part6_2-SCHEMATIC1-test.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 1 700m 700m
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\part6_2-SCHEMATIC1.net" 


.END
