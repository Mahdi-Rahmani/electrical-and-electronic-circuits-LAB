** Profile: "SCHEMATIC1-tes"  [ C:\USERS\M R\DESKTOP\AZ MADAR ELEC\6\S06\pishgozaresh\pish-SCHEMATIC1-tes.sim ] 

** Creating circuit file "pish-SCHEMATIC1-tes.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 0.1ms 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\pish-SCHEMATIC1.net" 


.END
