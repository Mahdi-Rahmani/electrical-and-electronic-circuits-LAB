** Profile: "SCHEMATIC1-test"  [ C:\USERS\M R\DESKTOP\AZ MADAR ELEC\s10\pish2\pish2-SCHEMATIC1-test.sim ] 

** Creating circuit file "pish2-SCHEMATIC1-test.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 3ms 0 3u 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\pish2-SCHEMATIC1.net" 


.END
