** Profile: "SCHEMATIC1-test"  [ C:\USERS\M R\DESKTOP\AZ MADAR ELEC\s10\pish7\pish6-SCHEMATIC1-test.sim ] 

** Creating circuit file "pish6-SCHEMATIC1-test.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 1000 0.001 30k
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\pish6-SCHEMATIC1.net" 


.END
