** Profile: "SCHEMATIC1-test2"  [ C:\USERS\M R\DESKTOP\AZ MADAR ELEC\elec project\q4\part4-SCHEMATIC1-test2.sim ] 

** Creating circuit file "part4-SCHEMATIC1-test2.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN PARAM a 10m 50m 5m 
+ LIN PARAM b 10m 50m 5m 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\part4-SCHEMATIC1.net" 


.END
