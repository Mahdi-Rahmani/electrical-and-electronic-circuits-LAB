** Profile: "SCHEMATIC1-te1"  [ C:\USERS\M R\DESKTOP\az madar elec\s07\azmayesh4\az4-SCHEMATIC1-te1.sim ] 

** Creating circuit file "az4-SCHEMATIC1-te1.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 1000 0.1 200k
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\az4-SCHEMATIC1.net" 


.END
