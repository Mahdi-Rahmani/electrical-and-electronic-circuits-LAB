** Profile: "SCHEMATIC1-test"  [ C:\USERS\M R\DESKTOP\AZ MADAR ELEC\6\S06\azmayesh 3\az3-SCHEMATIC1-test.sim ] 

** Creating circuit file "az3-SCHEMATIC1-test.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 0.06ms 0 
.STEP LIN PARAM a 10k 11k 0.2k 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\az3-SCHEMATIC1.net" 


.END
