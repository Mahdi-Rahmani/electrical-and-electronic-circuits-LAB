** Profile: "SCHEMATIC1-tes2"  [ C:\USERS\M R\DESKTOP\AZ MADAR ELEC\s09\az4\az4-SCHEMATIC1-tes2.sim ] 

** Creating circuit file "az4-SCHEMATIC1-tes2.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1ms 0 1u 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\az4-SCHEMATIC1.net" 


.END
