** Profile: "SCHEMATIC1-q4-simulat"  [ C:\USERS\M R\DESKTOP\AZ MADAR ELEC\pishgozaresh\q3\q4_pishgozaresh-SCHEMATIC1-q4-simulat.sim ] 

** Creating circuit file "q4_pishgozaresh-SCHEMATIC1-q4-simulat.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\q4_pishgozaresh-SCHEMATIC1.net" 


.END
