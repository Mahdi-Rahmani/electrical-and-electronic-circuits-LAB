** Profile: "SCHEMATIC1-tast"  [ C:\Users\M R\Desktop\az madar elec\6\s06\azmayesh 1\q1-SCHEMATIC1-tast.sim ] 

** Creating circuit file "q1-SCHEMATIC1-tast.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 0.2ms 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\q1-SCHEMATIC1.net" 


.END
