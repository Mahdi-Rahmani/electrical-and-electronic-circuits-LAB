** Profile: "SCHEMATIC1-az1"  [ C:\Users\M R\Desktop\az madar elec\se2\s02\s02-schematic1-az1.sim ] 

** Creating circuit file "s02-schematic1-az1.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN PARAM a 0 1 0.2 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\s02-SCHEMATIC1.net" 


.END
