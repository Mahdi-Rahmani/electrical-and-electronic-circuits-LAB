** Profile: "SCHEMATIC1-test"  [ C:\USERS\M R\DESKTOP\AZ MADAR ELEC\elec project\q5\part5-SCHEMATIC1-test.sim ] 

** Creating circuit file "part5-SCHEMATIC1-test.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 10000 1u 100k
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\part5-SCHEMATIC1.net" 


.END
