** Profile: "SCHEMATIC1-test2"  [ C:\Users\M R\Desktop\az madar elec\s03\pish gozaresh 2\soal4\part1\level1\q4-1-SCHEMATIC1-test2.sim ] 

** Creating circuit file "q4-1-SCHEMATIC1-test2.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1000ns 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\q4-1-SCHEMATIC1.net" 


.END
