** Profile: "SCHEMATIC1-test"  [ C:\Users\M R\Desktop\az madar elec\6\s06\azmayesh 5\az5-schematic1-test.sim ] 

** Creating circuit file "az5-schematic1-test.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 0.5ms 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\az5-SCHEMATIC1.net" 


.END
