** Profile: "SCHEMATIC1-test"  [ C:\Users\M R\Desktop\az madar elec\s05\part1\pish gozaresh2\q2-SCHEMATIC1-test.sim ] 

** Creating circuit file "q2-SCHEMATIC1-test.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 40ms 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\q2-SCHEMATIC1.net" 


.END
