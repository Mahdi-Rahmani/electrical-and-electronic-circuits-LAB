** Profile: "SCHEMATIC1-tets"  [ C:\USERS\M R\DESKTOP\AZ MADAR ELEC\ELEC PROJECT\Q6\SECOND STATE\I\in-SCHEMATIC1-tets.sim ] 

** Creating circuit file "in-SCHEMATIC1-tets.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 1 700m 700m
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\in-SCHEMATIC1.net" 


.END
