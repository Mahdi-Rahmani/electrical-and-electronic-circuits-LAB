** Profile: "SCHEMATIC1-dc"  [ C:\USERS\M R\DESKTOP\az madar elec\s07\pishGozaresh1\pish1-SCHEMATIC1-dc.sim ] 

** Creating circuit file "pish1-SCHEMATIC1-dc.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\pish1-SCHEMATIC1.net" 


.END
