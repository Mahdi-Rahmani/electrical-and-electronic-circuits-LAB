** Profile: "SCHEMATIC1-test1"  [ C:\Users\M R\Desktop\az madar elec\s05\part1\azmayesh1\q1-SCHEMATIC1-test1.sim ] 

** Creating circuit file "q1-SCHEMATIC1-test1.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 60ms 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\q1-SCHEMATIC1.net" 


.END
