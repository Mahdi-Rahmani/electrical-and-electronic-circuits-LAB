** Profile: "SCHEMATIC1-test"  [ C:\USERS\M R\DESKTOP\az madar elec\s07\pishgozaresh3\q3-SCHEMATIC1-test.sim ] 

** Creating circuit file "q3-SCHEMATIC1-test.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 10ms 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\q3-SCHEMATIC1.net" 


.END
