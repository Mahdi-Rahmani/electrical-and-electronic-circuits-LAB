** Profile: "SCHEMATIC1-pish1Sim"  [ C:\USERS\M R\DESKTOP\az madar elec\s07\pishGozaresh1\pish1-SCHEMATIC1-pish1Sim.sim ] 

** Creating circuit file "pish1-SCHEMATIC1-pish1Sim.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 1000 0.1 200k
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\pish1-SCHEMATIC1.net" 


.END
